// Qsys.v

// Generated using ACDS version 16.0 222

`timescale 1 ps / 1 ps
module Qsys (
		input  wire        bts_tmd_connect_state_external_connection_export, // bts_tmd_connect_state_external_connection.export
		output wire        buzzer_out_external_connection_export,            //            buzzer_out_external_connection.export
		output wire [1:0]  car_led_external_connection_export,               //               car_led_external_connection.export
		input  wire [11:0] car_voltage_data_external_connection_export,      //      car_voltage_data_external_connection.export
		input  wire        clk_clk,                                          //                                       clk.clk
		output wire        dc_motor_left_conduit_end_motor_p,                //                 dc_motor_left_conduit_end.motor_p
		output wire        dc_motor_left_conduit_end_motor_n,                //                                          .motor_n
		output wire        dc_motor_right_conduit_end_motor_p,               //                dc_motor_right_conduit_end.motor_p
		output wire        dc_motor_right_conduit_end_motor_n,               //                                          .motor_n
		output wire [7:0]  led_external_connection_export,                   //                   led_external_connection.export
		input  wire [1:0]  motor_measure_left_conduit_end_ab,                //            motor_measure_left_conduit_end.ab
		input  wire [1:0]  motor_measure_right_conduit_end_ab,               //           motor_measure_right_conduit_end.ab
		inout  wire        mpu_i2c_export_scl_pad_io,                        //                            mpu_i2c_export.scl_pad_io
		inout  wire        mpu_i2c_export_sda_pad_io,                        //                                          .sda_pad_io
		input  wire        mpu_int_external_connection_export,               //               mpu_int_external_connection.export
		input  wire        pmonitor_alert_external_connection_export,        //        pmonitor_alert_external_connection.export
		inout  wire        pwmonitor_i2c_export_scl_pad_io,                  //                      pwmonitor_i2c_export.scl_pad_io
		inout  wire        pwmonitor_i2c_export_sda_pad_io,                  //                                          .sda_pad_io
		input  wire        reset_reset_n,                                    //                                     reset.reset_n
		input  wire        sonic_distance_0_conduit_end_echo,                //              sonic_distance_0_conduit_end.echo
		output wire        sonic_distance_0_conduit_end_trigger,             //                                          .trigger
		input  wire        uart_bt_external_interface_RXD,                   //                uart_bt_external_interface.RXD
		output wire        uart_bt_external_interface_TXD                    //                                          .TXD
	);

	wire         pll_0_outclk0_clk;                                               // pll_0:outclk_0 -> [bts_tmd_connect_state:clk, buzzer_out:clk, car_led:clk, car_voltage_data:clk, dc_motor_left:clk, dc_motor_right:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, mm_clock_crossing_bridge_0:s0_clk, mm_interconnect_0:pll_0_outclk0_clk, motor_measure_left:clk, motor_measure_right:clk, mpu_int:clk, nios2_gen2_0:clk, onchip_memory2_0:clk, rst_controller_001:clk, rst_controller_002:clk, sysid_qsys:clock, timer_0:clk]
	wire         pll_0_outclk1_clk;                                               // pll_0:outclk_1 -> [mm_interconnect_0:pll_0_outclk1_clk, pmonitor_alert:clk, rst_controller_003:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                               // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                            // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                            // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [24:0] nios2_gen2_0_data_master_address;                                // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                             // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                   // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                                  // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                              // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                        // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                     // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [24:0] nios2_gen2_0_instruction_master_address;                         // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                            // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;          // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;       // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_uart_bt_avalon_rs232_slave_chipselect;         // mm_interconnect_0:uart_bt_avalon_rs232_slave_chipselect -> uart_bt:chipselect
	wire  [31:0] mm_interconnect_0_uart_bt_avalon_rs232_slave_readdata;           // uart_bt:readdata -> mm_interconnect_0:uart_bt_avalon_rs232_slave_readdata
	wire   [0:0] mm_interconnect_0_uart_bt_avalon_rs232_slave_address;            // mm_interconnect_0:uart_bt_avalon_rs232_slave_address -> uart_bt:address
	wire         mm_interconnect_0_uart_bt_avalon_rs232_slave_read;               // mm_interconnect_0:uart_bt_avalon_rs232_slave_read -> uart_bt:read
	wire   [3:0] mm_interconnect_0_uart_bt_avalon_rs232_slave_byteenable;         // mm_interconnect_0:uart_bt_avalon_rs232_slave_byteenable -> uart_bt:byteenable
	wire         mm_interconnect_0_uart_bt_avalon_rs232_slave_write;              // mm_interconnect_0:uart_bt_avalon_rs232_slave_write -> uart_bt:write
	wire  [31:0] mm_interconnect_0_uart_bt_avalon_rs232_slave_writedata;          // mm_interconnect_0:uart_bt_avalon_rs232_slave_writedata -> uart_bt:writedata
	wire         mm_interconnect_0_dc_motor_left_avalon_slave_chipselect;         // mm_interconnect_0:dc_motor_left_avalon_slave_chipselect -> dc_motor_left:s_cs
	wire  [31:0] mm_interconnect_0_dc_motor_left_avalon_slave_readdata;           // dc_motor_left:s_readdata -> mm_interconnect_0:dc_motor_left_avalon_slave_readdata
	wire   [1:0] mm_interconnect_0_dc_motor_left_avalon_slave_address;            // mm_interconnect_0:dc_motor_left_avalon_slave_address -> dc_motor_left:s_address
	wire         mm_interconnect_0_dc_motor_left_avalon_slave_read;               // mm_interconnect_0:dc_motor_left_avalon_slave_read -> dc_motor_left:s_read
	wire         mm_interconnect_0_dc_motor_left_avalon_slave_write;              // mm_interconnect_0:dc_motor_left_avalon_slave_write -> dc_motor_left:s_write
	wire  [31:0] mm_interconnect_0_dc_motor_left_avalon_slave_writedata;          // mm_interconnect_0:dc_motor_left_avalon_slave_writedata -> dc_motor_left:s_writedata
	wire         mm_interconnect_0_dc_motor_right_avalon_slave_chipselect;        // mm_interconnect_0:dc_motor_right_avalon_slave_chipselect -> dc_motor_right:s_cs
	wire  [31:0] mm_interconnect_0_dc_motor_right_avalon_slave_readdata;          // dc_motor_right:s_readdata -> mm_interconnect_0:dc_motor_right_avalon_slave_readdata
	wire   [1:0] mm_interconnect_0_dc_motor_right_avalon_slave_address;           // mm_interconnect_0:dc_motor_right_avalon_slave_address -> dc_motor_right:s_address
	wire         mm_interconnect_0_dc_motor_right_avalon_slave_read;              // mm_interconnect_0:dc_motor_right_avalon_slave_read -> dc_motor_right:s_read
	wire         mm_interconnect_0_dc_motor_right_avalon_slave_write;             // mm_interconnect_0:dc_motor_right_avalon_slave_write -> dc_motor_right:s_write
	wire  [31:0] mm_interconnect_0_dc_motor_right_avalon_slave_writedata;         // mm_interconnect_0:dc_motor_right_avalon_slave_writedata -> dc_motor_right:s_writedata
	wire         mm_interconnect_0_motor_measure_left_avalon_slave_0_chipselect;  // mm_interconnect_0:motor_measure_left_avalon_slave_0_chipselect -> motor_measure_left:s_cs
	wire  [31:0] mm_interconnect_0_motor_measure_left_avalon_slave_0_readdata;    // motor_measure_left:s_readdata -> mm_interconnect_0:motor_measure_left_avalon_slave_0_readdata
	wire   [2:0] mm_interconnect_0_motor_measure_left_avalon_slave_0_address;     // mm_interconnect_0:motor_measure_left_avalon_slave_0_address -> motor_measure_left:s_address
	wire         mm_interconnect_0_motor_measure_left_avalon_slave_0_read;        // mm_interconnect_0:motor_measure_left_avalon_slave_0_read -> motor_measure_left:s_read
	wire         mm_interconnect_0_motor_measure_left_avalon_slave_0_write;       // mm_interconnect_0:motor_measure_left_avalon_slave_0_write -> motor_measure_left:s_write
	wire  [31:0] mm_interconnect_0_motor_measure_left_avalon_slave_0_writedata;   // mm_interconnect_0:motor_measure_left_avalon_slave_0_writedata -> motor_measure_left:s_writedata
	wire         mm_interconnect_0_motor_measure_right_avalon_slave_0_chipselect; // mm_interconnect_0:motor_measure_right_avalon_slave_0_chipselect -> motor_measure_right:s_cs
	wire  [31:0] mm_interconnect_0_motor_measure_right_avalon_slave_0_readdata;   // motor_measure_right:s_readdata -> mm_interconnect_0:motor_measure_right_avalon_slave_0_readdata
	wire   [2:0] mm_interconnect_0_motor_measure_right_avalon_slave_0_address;    // mm_interconnect_0:motor_measure_right_avalon_slave_0_address -> motor_measure_right:s_address
	wire         mm_interconnect_0_motor_measure_right_avalon_slave_0_read;       // mm_interconnect_0:motor_measure_right_avalon_slave_0_read -> motor_measure_right:s_read
	wire         mm_interconnect_0_motor_measure_right_avalon_slave_0_write;      // mm_interconnect_0:motor_measure_right_avalon_slave_0_write -> motor_measure_right:s_write
	wire  [31:0] mm_interconnect_0_motor_measure_right_avalon_slave_0_writedata;  // mm_interconnect_0:motor_measure_right_avalon_slave_0_writedata -> motor_measure_right:s_writedata
	wire         mm_interconnect_0_mpu_i2c_avalon_slave_0_chipselect;             // mm_interconnect_0:mpu_i2c_avalon_slave_0_chipselect -> mpu_i2c:wb_stb_i
	wire   [7:0] mm_interconnect_0_mpu_i2c_avalon_slave_0_readdata;               // mpu_i2c:wb_dat_o -> mm_interconnect_0:mpu_i2c_avalon_slave_0_readdata
	wire         mm_interconnect_0_mpu_i2c_avalon_slave_0_waitrequest;            // mpu_i2c:wb_ack_o -> mm_interconnect_0:mpu_i2c_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_mpu_i2c_avalon_slave_0_address;                // mm_interconnect_0:mpu_i2c_avalon_slave_0_address -> mpu_i2c:wb_adr_i
	wire         mm_interconnect_0_mpu_i2c_avalon_slave_0_write;                  // mm_interconnect_0:mpu_i2c_avalon_slave_0_write -> mpu_i2c:wb_we_i
	wire   [7:0] mm_interconnect_0_mpu_i2c_avalon_slave_0_writedata;              // mm_interconnect_0:mpu_i2c_avalon_slave_0_writedata -> mpu_i2c:wb_dat_i
	wire         mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_chipselect;       // mm_interconnect_0:pwmonitor_i2c_avalon_slave_0_chipselect -> pwmonitor_i2c:wb_stb_i
	wire   [7:0] mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_readdata;         // pwmonitor_i2c:wb_dat_o -> mm_interconnect_0:pwmonitor_i2c_avalon_slave_0_readdata
	wire         mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_waitrequest;      // pwmonitor_i2c:wb_ack_o -> mm_interconnect_0:pwmonitor_i2c_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_address;          // mm_interconnect_0:pwmonitor_i2c_avalon_slave_0_address -> pwmonitor_i2c:wb_adr_i
	wire         mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_write;            // mm_interconnect_0:pwmonitor_i2c_avalon_slave_0_write -> pwmonitor_i2c:wb_we_i
	wire   [7:0] mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_writedata;        // mm_interconnect_0:pwmonitor_i2c_avalon_slave_0_writedata -> pwmonitor_i2c:wb_dat_i
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;             // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;              // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;         // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;      // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;             // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata;        // mm_clock_crossing_bridge_0:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest;     // mm_clock_crossing_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess;     // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_debugaccess -> mm_clock_crossing_bridge_0:s0_debugaccess
	wire   [4:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address;         // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_address -> mm_clock_crossing_bridge_0:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read;            // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_read -> mm_clock_crossing_bridge_0:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable;      // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_byteenable -> mm_clock_crossing_bridge_0:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid;   // mm_clock_crossing_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write;           // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_write -> mm_clock_crossing_bridge_0:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata;       // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_writedata -> mm_clock_crossing_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount;      // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_burstcount -> mm_clock_crossing_bridge_0:s0_burstcount
	wire         mm_interconnect_0_buzzer_out_s1_chipselect;                      // mm_interconnect_0:buzzer_out_s1_chipselect -> buzzer_out:chipselect
	wire  [31:0] mm_interconnect_0_buzzer_out_s1_readdata;                        // buzzer_out:readdata -> mm_interconnect_0:buzzer_out_s1_readdata
	wire   [1:0] mm_interconnect_0_buzzer_out_s1_address;                         // mm_interconnect_0:buzzer_out_s1_address -> buzzer_out:address
	wire         mm_interconnect_0_buzzer_out_s1_write;                           // mm_interconnect_0:buzzer_out_s1_write -> buzzer_out:write_n
	wire  [31:0] mm_interconnect_0_buzzer_out_s1_writedata;                       // mm_interconnect_0:buzzer_out_s1_writedata -> buzzer_out:writedata
	wire  [31:0] mm_interconnect_0_car_voltage_data_s1_readdata;                  // car_voltage_data:readdata -> mm_interconnect_0:car_voltage_data_s1_readdata
	wire   [1:0] mm_interconnect_0_car_voltage_data_s1_address;                   // mm_interconnect_0:car_voltage_data_s1_address -> car_voltage_data:address
	wire         mm_interconnect_0_car_led_s1_chipselect;                         // mm_interconnect_0:car_led_s1_chipselect -> car_led:chipselect
	wire  [31:0] mm_interconnect_0_car_led_s1_readdata;                           // car_led:readdata -> mm_interconnect_0:car_led_s1_readdata
	wire   [1:0] mm_interconnect_0_car_led_s1_address;                            // mm_interconnect_0:car_led_s1_address -> car_led:address
	wire         mm_interconnect_0_car_led_s1_write;                              // mm_interconnect_0:car_led_s1_write -> car_led:write_n
	wire  [31:0] mm_interconnect_0_car_led_s1_writedata;                          // mm_interconnect_0:car_led_s1_writedata -> car_led:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                         // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                           // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                            // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                              // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                          // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire  [31:0] mm_interconnect_0_bts_tmd_connect_state_s1_readdata;             // bts_tmd_connect_state:readdata -> mm_interconnect_0:bts_tmd_connect_state_s1_readdata
	wire   [1:0] mm_interconnect_0_bts_tmd_connect_state_s1_address;              // mm_interconnect_0:bts_tmd_connect_state_s1_address -> bts_tmd_connect_state:address
	wire         mm_interconnect_0_mpu_int_s1_chipselect;                         // mm_interconnect_0:mpu_int_s1_chipselect -> mpu_int:chipselect
	wire  [31:0] mm_interconnect_0_mpu_int_s1_readdata;                           // mpu_int:readdata -> mm_interconnect_0:mpu_int_s1_readdata
	wire   [1:0] mm_interconnect_0_mpu_int_s1_address;                            // mm_interconnect_0:mpu_int_s1_address -> mpu_int:address
	wire         mm_interconnect_0_mpu_int_s1_write;                              // mm_interconnect_0:mpu_int_s1_write -> mpu_int:write_n
	wire  [31:0] mm_interconnect_0_mpu_int_s1_writedata;                          // mm_interconnect_0:mpu_int_s1_writedata -> mpu_int:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                  // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_address;                   // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                     // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                 // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                     // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_pmonitor_alert_s1_readdata;                    // pmonitor_alert:readdata -> mm_interconnect_0:pmonitor_alert_s1_readdata
	wire   [1:0] mm_interconnect_0_pmonitor_alert_s1_address;                     // mm_interconnect_0:pmonitor_alert_s1_address -> pmonitor_alert:address
	wire         mm_clock_crossing_bridge_0_m0_waitrequest;                       // mm_interconnect_1:mm_clock_crossing_bridge_0_m0_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_0_m0_readdata;                          // mm_interconnect_1:mm_clock_crossing_bridge_0_m0_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	wire         mm_clock_crossing_bridge_0_m0_debugaccess;                       // mm_clock_crossing_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_debugaccess
	wire   [4:0] mm_clock_crossing_bridge_0_m0_address;                           // mm_clock_crossing_bridge_0:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_address
	wire         mm_clock_crossing_bridge_0_m0_read;                              // mm_clock_crossing_bridge_0:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_read
	wire   [3:0] mm_clock_crossing_bridge_0_m0_byteenable;                        // mm_clock_crossing_bridge_0:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_byteenable
	wire         mm_clock_crossing_bridge_0_m0_readdatavalid;                     // mm_interconnect_1:mm_clock_crossing_bridge_0_m0_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_0_m0_writedata;                         // mm_clock_crossing_bridge_0:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_writedata
	wire         mm_clock_crossing_bridge_0_m0_write;                             // mm_clock_crossing_bridge_0:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_write
	wire   [0:0] mm_clock_crossing_bridge_0_m0_burstcount;                        // mm_clock_crossing_bridge_0:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_burstcount
	wire         mm_interconnect_1_sonic_distance_0_avalon_slave_0_chipselect;    // mm_interconnect_1:sonic_distance_0_avalon_slave_0_chipselect -> sonic_distance_0:av_mm_cs
	wire  [31:0] mm_interconnect_1_sonic_distance_0_avalon_slave_0_readdata;      // sonic_distance_0:av_mm_readdata -> mm_interconnect_1:sonic_distance_0_avalon_slave_0_readdata
	wire   [0:0] mm_interconnect_1_sonic_distance_0_avalon_slave_0_address;       // mm_interconnect_1:sonic_distance_0_avalon_slave_0_address -> sonic_distance_0:av_mm_address
	wire         mm_interconnect_1_sonic_distance_0_avalon_slave_0_read;          // mm_interconnect_1:sonic_distance_0_avalon_slave_0_read -> sonic_distance_0:av_mm_read
	wire         mm_interconnect_1_led_s1_chipselect;                             // mm_interconnect_1:LED_s1_chipselect -> LED:chipselect
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                               // LED:readdata -> mm_interconnect_1:LED_s1_readdata
	wire   [1:0] mm_interconnect_1_led_s1_address;                                // mm_interconnect_1:LED_s1_address -> LED:address
	wire         mm_interconnect_1_led_s1_write;                                  // mm_interconnect_1:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                              // mm_interconnect_1:LED_s1_writedata -> LED:writedata
	wire         irq_mapper_receiver2_irq;                                        // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                        // timer_0:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                        // mpu_int:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                            // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         irq_mapper_receiver0_irq;                                        // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                   // uart_bt:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                        // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                               // pwmonitor_i2c:wb_inta_o -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [LED:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_clock_crossing_bridge_0:m0_reset, mm_interconnect_0:uart_bt_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset, mpu_i2c:wb_rst_i, pwmonitor_i2c:wb_rst_i, sonic_distance_0:av_mm_rst, uart_bt:reset]
	wire         rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [bts_tmd_connect_state:reset_n, buzzer_out:reset_n, car_led:reset_n, car_voltage_data:reset_n, dc_motor_left:reset_n, dc_motor_right:reset_n, jtag_uart:rst_n, mm_clock_crossing_bridge_0:s0_reset, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, motor_measure_left:reset_n, motor_measure_right:reset_n, mpu_int:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sysid_qsys:reset_n, timer_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                          // rst_controller_001:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                              // rst_controller_002:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator_001:in_reset]
	wire         rst_controller_002_reset_out_reset_req;                          // rst_controller_002:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                          // nios2_gen2_0:debug_reset_request -> rst_controller_002:reset_in1
	wire         rst_controller_003_reset_out_reset;                              // rst_controller_003:reset_out -> [mm_interconnect_0:pmonitor_alert_reset_reset_bridge_in_reset_reset, pmonitor_alert:reset_n]

	Qsys_LED led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	Qsys_bts_tmd_connect_state bts_tmd_connect_state (
		.clk      (pll_0_outclk0_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_bts_tmd_connect_state_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_bts_tmd_connect_state_s1_readdata), //                    .readdata
		.in_port  (bts_tmd_connect_state_external_connection_export)     // external_connection.export
	);

	Qsys_buzzer_out buzzer_out (
		.clk        (pll_0_outclk0_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_buzzer_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buzzer_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buzzer_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buzzer_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buzzer_out_s1_readdata),   //                    .readdata
		.out_port   (buzzer_out_external_connection_export)       // external_connection.export
	);

	Qsys_car_led car_led (
		.clk        (pll_0_outclk0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_car_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_car_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_car_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_car_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_car_led_s1_readdata),   //                    .readdata
		.out_port   (car_led_external_connection_export)       // external_connection.export
	);

	Qsys_car_voltage_data car_voltage_data (
		.clk      (pll_0_outclk0_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_car_voltage_data_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_car_voltage_data_s1_readdata), //                    .readdata
		.in_port  (car_voltage_data_external_connection_export)     // external_connection.export
	);

	Qsys_dc_motor_left dc_motor_left (
		.clk         (pll_0_outclk0_clk),                                       //        clock.clk
		.reset_n     (~rst_controller_001_reset_out_reset),                     //        reset.reset_n
		.s_cs        (mm_interconnect_0_dc_motor_left_avalon_slave_chipselect), // avalon_slave.chipselect
		.s_address   (mm_interconnect_0_dc_motor_left_avalon_slave_address),    //             .address
		.s_write     (mm_interconnect_0_dc_motor_left_avalon_slave_write),      //             .write
		.s_writedata (mm_interconnect_0_dc_motor_left_avalon_slave_writedata),  //             .writedata
		.s_read      (mm_interconnect_0_dc_motor_left_avalon_slave_read),       //             .read
		.s_readdata  (mm_interconnect_0_dc_motor_left_avalon_slave_readdata),   //             .readdata
		.DC_MOTOR_P  (dc_motor_left_conduit_end_motor_p),                       //  conduit_end.motor_p
		.DC_MOTOR_N  (dc_motor_left_conduit_end_motor_n)                        //             .motor_n
	);

	Qsys_dc_motor_left dc_motor_right (
		.clk         (pll_0_outclk0_clk),                                        //        clock.clk
		.reset_n     (~rst_controller_001_reset_out_reset),                      //        reset.reset_n
		.s_cs        (mm_interconnect_0_dc_motor_right_avalon_slave_chipselect), // avalon_slave.chipselect
		.s_address   (mm_interconnect_0_dc_motor_right_avalon_slave_address),    //             .address
		.s_write     (mm_interconnect_0_dc_motor_right_avalon_slave_write),      //             .write
		.s_writedata (mm_interconnect_0_dc_motor_right_avalon_slave_writedata),  //             .writedata
		.s_read      (mm_interconnect_0_dc_motor_right_avalon_slave_read),       //             .read
		.s_readdata  (mm_interconnect_0_dc_motor_right_avalon_slave_readdata),   //             .readdata
		.DC_MOTOR_P  (dc_motor_right_conduit_end_motor_p),                       //  conduit_end.motor_p
		.DC_MOTOR_N  (dc_motor_right_conduit_end_motor_n)                        //             .motor_n
	);

	Qsys_jtag_uart jtag_uart (
		.clk            (pll_0_outclk0_clk),                                         //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (5),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (16),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_0 (
		.m0_clk           (clk_clk),                                                       //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                                // m0_reset.reset
		.s0_clk           (pll_0_outclk0_clk),                                             //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                            // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_0_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_0_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_0_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_0_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_0_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_0_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_0_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_0_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_0_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_0_m0_debugaccess)                      //         .debugaccess
	);

	Qsys_motor_measure_left motor_measure_left (
		.s_cs        (mm_interconnect_0_motor_measure_left_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.s_write     (mm_interconnect_0_motor_measure_left_avalon_slave_0_write),      //               .write
		.s_read      (mm_interconnect_0_motor_measure_left_avalon_slave_0_read),       //               .read
		.s_address   (mm_interconnect_0_motor_measure_left_avalon_slave_0_address),    //               .address
		.s_writedata (mm_interconnect_0_motor_measure_left_avalon_slave_0_writedata),  //               .writedata
		.s_readdata  (mm_interconnect_0_motor_measure_left_avalon_slave_0_readdata),   //               .readdata
		.clk         (pll_0_outclk0_clk),                                              //          clock.clk
		.reset_n     (~rst_controller_001_reset_out_reset),                            //          reset.reset_n
		.phase_AB    (motor_measure_left_conduit_end_ab)                               //    conduit_end.ab
	);

	Qsys_motor_measure_left motor_measure_right (
		.s_cs        (mm_interconnect_0_motor_measure_right_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.s_write     (mm_interconnect_0_motor_measure_right_avalon_slave_0_write),      //               .write
		.s_read      (mm_interconnect_0_motor_measure_right_avalon_slave_0_read),       //               .read
		.s_address   (mm_interconnect_0_motor_measure_right_avalon_slave_0_address),    //               .address
		.s_writedata (mm_interconnect_0_motor_measure_right_avalon_slave_0_writedata),  //               .writedata
		.s_readdata  (mm_interconnect_0_motor_measure_right_avalon_slave_0_readdata),   //               .readdata
		.clk         (pll_0_outclk0_clk),                                               //          clock.clk
		.reset_n     (~rst_controller_001_reset_out_reset),                             //          reset.reset_n
		.phase_AB    (motor_measure_right_conduit_end_ab)                               //    conduit_end.ab
	);

	i2c_opencores mpu_i2c (
		.wb_clk_i   (clk_clk),                                              //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                       //      clock_reset.reset
		.scl_pad_io (mpu_i2c_export_scl_pad_io),                            //           export.export
		.sda_pad_io (mpu_i2c_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_mpu_i2c_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_mpu_i2c_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_mpu_i2c_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_mpu_i2c_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_mpu_i2c_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_mpu_i2c_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  ()                                                      // interrupt_sender.irq
	);

	Qsys_mpu_int mpu_int (
		.clk        (pll_0_outclk0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_mpu_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_mpu_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_mpu_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_mpu_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_mpu_int_s1_readdata),   //                    .readdata
		.in_port    (mpu_int_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                 //                 irq.irq
	);

	Qsys_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (pll_0_outclk0_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	Qsys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (pll_0_outclk0_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)            //       .reset_req
	);

	Qsys_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk), // outclk1.clk
		.locked   ()                   //  locked.export
	);

	Qsys_pmonitor_alert pmonitor_alert (
		.clk      (pll_0_outclk1_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pmonitor_alert_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pmonitor_alert_s1_readdata), //                    .readdata
		.in_port  (pmonitor_alert_external_connection_export)     // external_connection.export
	);

	i2c_opencores pwmonitor_i2c (
		.wb_clk_i   (clk_clk),                                                    //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                             //      clock_reset.reset
		.scl_pad_io (pwmonitor_i2c_export_scl_pad_io),                            //           export.export
		.sda_pad_io (pwmonitor_i2c_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_synchronizer_001_receiver_irq)                           // interrupt_sender.irq
	);

	Qsys_sonic_distance_0 sonic_distance_0 (
		.av_mm_cs       (mm_interconnect_1_sonic_distance_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.av_mm_address  (mm_interconnect_1_sonic_distance_0_avalon_slave_0_address),    //               .address
		.av_mm_read     (mm_interconnect_1_sonic_distance_0_avalon_slave_0_read),       //               .read
		.av_mm_readdata (mm_interconnect_1_sonic_distance_0_avalon_slave_0_readdata),   //               .readdata
		.av_mm_clk      (clk_clk),                                                      //     clock_sink.clk
		.av_mm_rst      (~rst_controller_reset_out_reset),                              //     reset_sink.reset_n
		.sonic_echo     (sonic_distance_0_conduit_end_echo),                            //    conduit_end.echo
		.sonic_trigger  (sonic_distance_0_conduit_end_trigger)                          //               .trigger
	);

	Qsys_sysid_qsys sysid_qsys (
		.clock    (pll_0_outclk0_clk),                                   //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	Qsys_timer_0 timer_0 (
		.clk        (pll_0_outclk0_clk),                       //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	Qsys_uart_bt uart_bt (
		.clk        (clk_clk),                                                 //                clk.clk
		.reset      (rst_controller_reset_out_reset),                          //              reset.reset
		.address    (mm_interconnect_0_uart_bt_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_uart_bt_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_uart_bt_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_uart_bt_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_uart_bt_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_uart_bt_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_uart_bt_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (irq_synchronizer_receiver_irq),                           //          interrupt.irq
		.UART_RXD   (uart_bt_external_interface_RXD),                          // external_interface.export
		.UART_TXD   (uart_bt_external_interface_TXD)                           //                   .export
	);

	Qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                         //                                  clk_0_clk.clk
		.pll_0_outclk0_clk                                (pll_0_outclk0_clk),                                               //                              pll_0_outclk0.clk
		.pll_0_outclk1_clk                                (pll_0_outclk1_clk),                                               //                              pll_0_outclk1.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                              //      jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset   (rst_controller_002_reset_out_reset),                              //   nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.pmonitor_alert_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                              // pmonitor_alert_reset_reset_bridge_in_reset.reset
		.uart_bt_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                                  //        uart_bt_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                 (nios2_gen2_0_data_master_address),                                //                   nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest             (nios2_gen2_0_data_master_waitrequest),                            //                                           .waitrequest
		.nios2_gen2_0_data_master_byteenable              (nios2_gen2_0_data_master_byteenable),                             //                                           .byteenable
		.nios2_gen2_0_data_master_read                    (nios2_gen2_0_data_master_read),                                   //                                           .read
		.nios2_gen2_0_data_master_readdata                (nios2_gen2_0_data_master_readdata),                               //                                           .readdata
		.nios2_gen2_0_data_master_readdatavalid           (nios2_gen2_0_data_master_readdatavalid),                          //                                           .readdatavalid
		.nios2_gen2_0_data_master_write                   (nios2_gen2_0_data_master_write),                                  //                                           .write
		.nios2_gen2_0_data_master_writedata               (nios2_gen2_0_data_master_writedata),                              //                                           .writedata
		.nios2_gen2_0_data_master_debugaccess             (nios2_gen2_0_data_master_debugaccess),                            //                                           .debugaccess
		.nios2_gen2_0_instruction_master_address          (nios2_gen2_0_instruction_master_address),                         //            nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest      (nios2_gen2_0_instruction_master_waitrequest),                     //                                           .waitrequest
		.nios2_gen2_0_instruction_master_read             (nios2_gen2_0_instruction_master_read),                            //                                           .read
		.nios2_gen2_0_instruction_master_readdata         (nios2_gen2_0_instruction_master_readdata),                        //                                           .readdata
		.nios2_gen2_0_instruction_master_readdatavalid    (nios2_gen2_0_instruction_master_readdatavalid),                   //                                           .readdatavalid
		.bts_tmd_connect_state_s1_address                 (mm_interconnect_0_bts_tmd_connect_state_s1_address),              //                   bts_tmd_connect_state_s1.address
		.bts_tmd_connect_state_s1_readdata                (mm_interconnect_0_bts_tmd_connect_state_s1_readdata),             //                                           .readdata
		.buzzer_out_s1_address                            (mm_interconnect_0_buzzer_out_s1_address),                         //                              buzzer_out_s1.address
		.buzzer_out_s1_write                              (mm_interconnect_0_buzzer_out_s1_write),                           //                                           .write
		.buzzer_out_s1_readdata                           (mm_interconnect_0_buzzer_out_s1_readdata),                        //                                           .readdata
		.buzzer_out_s1_writedata                          (mm_interconnect_0_buzzer_out_s1_writedata),                       //                                           .writedata
		.buzzer_out_s1_chipselect                         (mm_interconnect_0_buzzer_out_s1_chipselect),                      //                                           .chipselect
		.car_led_s1_address                               (mm_interconnect_0_car_led_s1_address),                            //                                 car_led_s1.address
		.car_led_s1_write                                 (mm_interconnect_0_car_led_s1_write),                              //                                           .write
		.car_led_s1_readdata                              (mm_interconnect_0_car_led_s1_readdata),                           //                                           .readdata
		.car_led_s1_writedata                             (mm_interconnect_0_car_led_s1_writedata),                          //                                           .writedata
		.car_led_s1_chipselect                            (mm_interconnect_0_car_led_s1_chipselect),                         //                                           .chipselect
		.car_voltage_data_s1_address                      (mm_interconnect_0_car_voltage_data_s1_address),                   //                        car_voltage_data_s1.address
		.car_voltage_data_s1_readdata                     (mm_interconnect_0_car_voltage_data_s1_readdata),                  //                                           .readdata
		.dc_motor_left_avalon_slave_address               (mm_interconnect_0_dc_motor_left_avalon_slave_address),            //                 dc_motor_left_avalon_slave.address
		.dc_motor_left_avalon_slave_write                 (mm_interconnect_0_dc_motor_left_avalon_slave_write),              //                                           .write
		.dc_motor_left_avalon_slave_read                  (mm_interconnect_0_dc_motor_left_avalon_slave_read),               //                                           .read
		.dc_motor_left_avalon_slave_readdata              (mm_interconnect_0_dc_motor_left_avalon_slave_readdata),           //                                           .readdata
		.dc_motor_left_avalon_slave_writedata             (mm_interconnect_0_dc_motor_left_avalon_slave_writedata),          //                                           .writedata
		.dc_motor_left_avalon_slave_chipselect            (mm_interconnect_0_dc_motor_left_avalon_slave_chipselect),         //                                           .chipselect
		.dc_motor_right_avalon_slave_address              (mm_interconnect_0_dc_motor_right_avalon_slave_address),           //                dc_motor_right_avalon_slave.address
		.dc_motor_right_avalon_slave_write                (mm_interconnect_0_dc_motor_right_avalon_slave_write),             //                                           .write
		.dc_motor_right_avalon_slave_read                 (mm_interconnect_0_dc_motor_right_avalon_slave_read),              //                                           .read
		.dc_motor_right_avalon_slave_readdata             (mm_interconnect_0_dc_motor_right_avalon_slave_readdata),          //                                           .readdata
		.dc_motor_right_avalon_slave_writedata            (mm_interconnect_0_dc_motor_right_avalon_slave_writedata),         //                                           .writedata
		.dc_motor_right_avalon_slave_chipselect           (mm_interconnect_0_dc_motor_right_avalon_slave_chipselect),        //                                           .chipselect
		.jtag_uart_avalon_jtag_slave_address              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),           //                jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),             //                                           .write
		.jtag_uart_avalon_jtag_slave_read                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),              //                                           .read
		.jtag_uart_avalon_jtag_slave_readdata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),          //                                           .readdata
		.jtag_uart_avalon_jtag_slave_writedata            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),         //                                           .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),       //                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),        //                                           .chipselect
		.mm_clock_crossing_bridge_0_s0_address            (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address),         //              mm_clock_crossing_bridge_0_s0.address
		.mm_clock_crossing_bridge_0_s0_write              (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write),           //                                           .write
		.mm_clock_crossing_bridge_0_s0_read               (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read),            //                                           .read
		.mm_clock_crossing_bridge_0_s0_readdata           (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata),        //                                           .readdata
		.mm_clock_crossing_bridge_0_s0_writedata          (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata),       //                                           .writedata
		.mm_clock_crossing_bridge_0_s0_burstcount         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount),      //                                           .burstcount
		.mm_clock_crossing_bridge_0_s0_byteenable         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable),      //                                           .byteenable
		.mm_clock_crossing_bridge_0_s0_readdatavalid      (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid),   //                                           .readdatavalid
		.mm_clock_crossing_bridge_0_s0_waitrequest        (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest),     //                                           .waitrequest
		.mm_clock_crossing_bridge_0_s0_debugaccess        (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess),     //                                           .debugaccess
		.motor_measure_left_avalon_slave_0_address        (mm_interconnect_0_motor_measure_left_avalon_slave_0_address),     //          motor_measure_left_avalon_slave_0.address
		.motor_measure_left_avalon_slave_0_write          (mm_interconnect_0_motor_measure_left_avalon_slave_0_write),       //                                           .write
		.motor_measure_left_avalon_slave_0_read           (mm_interconnect_0_motor_measure_left_avalon_slave_0_read),        //                                           .read
		.motor_measure_left_avalon_slave_0_readdata       (mm_interconnect_0_motor_measure_left_avalon_slave_0_readdata),    //                                           .readdata
		.motor_measure_left_avalon_slave_0_writedata      (mm_interconnect_0_motor_measure_left_avalon_slave_0_writedata),   //                                           .writedata
		.motor_measure_left_avalon_slave_0_chipselect     (mm_interconnect_0_motor_measure_left_avalon_slave_0_chipselect),  //                                           .chipselect
		.motor_measure_right_avalon_slave_0_address       (mm_interconnect_0_motor_measure_right_avalon_slave_0_address),    //         motor_measure_right_avalon_slave_0.address
		.motor_measure_right_avalon_slave_0_write         (mm_interconnect_0_motor_measure_right_avalon_slave_0_write),      //                                           .write
		.motor_measure_right_avalon_slave_0_read          (mm_interconnect_0_motor_measure_right_avalon_slave_0_read),       //                                           .read
		.motor_measure_right_avalon_slave_0_readdata      (mm_interconnect_0_motor_measure_right_avalon_slave_0_readdata),   //                                           .readdata
		.motor_measure_right_avalon_slave_0_writedata     (mm_interconnect_0_motor_measure_right_avalon_slave_0_writedata),  //                                           .writedata
		.motor_measure_right_avalon_slave_0_chipselect    (mm_interconnect_0_motor_measure_right_avalon_slave_0_chipselect), //                                           .chipselect
		.mpu_i2c_avalon_slave_0_address                   (mm_interconnect_0_mpu_i2c_avalon_slave_0_address),                //                     mpu_i2c_avalon_slave_0.address
		.mpu_i2c_avalon_slave_0_write                     (mm_interconnect_0_mpu_i2c_avalon_slave_0_write),                  //                                           .write
		.mpu_i2c_avalon_slave_0_readdata                  (mm_interconnect_0_mpu_i2c_avalon_slave_0_readdata),               //                                           .readdata
		.mpu_i2c_avalon_slave_0_writedata                 (mm_interconnect_0_mpu_i2c_avalon_slave_0_writedata),              //                                           .writedata
		.mpu_i2c_avalon_slave_0_waitrequest               (~mm_interconnect_0_mpu_i2c_avalon_slave_0_waitrequest),           //                                           .waitrequest
		.mpu_i2c_avalon_slave_0_chipselect                (mm_interconnect_0_mpu_i2c_avalon_slave_0_chipselect),             //                                           .chipselect
		.mpu_int_s1_address                               (mm_interconnect_0_mpu_int_s1_address),                            //                                 mpu_int_s1.address
		.mpu_int_s1_write                                 (mm_interconnect_0_mpu_int_s1_write),                              //                                           .write
		.mpu_int_s1_readdata                              (mm_interconnect_0_mpu_int_s1_readdata),                           //                                           .readdata
		.mpu_int_s1_writedata                             (mm_interconnect_0_mpu_int_s1_writedata),                          //                                           .writedata
		.mpu_int_s1_chipselect                            (mm_interconnect_0_mpu_int_s1_chipselect),                         //                                           .chipselect
		.nios2_gen2_0_debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),          //               nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),            //                                           .write
		.nios2_gen2_0_debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),             //                                           .read
		.nios2_gen2_0_debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),         //                                           .readdata
		.nios2_gen2_0_debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),        //                                           .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),       //                                           .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),      //                                           .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),      //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                   //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                     //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),                  //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),                 //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                     //                                           .clken
		.pmonitor_alert_s1_address                        (mm_interconnect_0_pmonitor_alert_s1_address),                     //                          pmonitor_alert_s1.address
		.pmonitor_alert_s1_readdata                       (mm_interconnect_0_pmonitor_alert_s1_readdata),                    //                                           .readdata
		.pwmonitor_i2c_avalon_slave_0_address             (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_address),          //               pwmonitor_i2c_avalon_slave_0.address
		.pwmonitor_i2c_avalon_slave_0_write               (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_write),            //                                           .write
		.pwmonitor_i2c_avalon_slave_0_readdata            (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_readdata),         //                                           .readdata
		.pwmonitor_i2c_avalon_slave_0_writedata           (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_writedata),        //                                           .writedata
		.pwmonitor_i2c_avalon_slave_0_waitrequest         (~mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_waitrequest),     //                                           .waitrequest
		.pwmonitor_i2c_avalon_slave_0_chipselect          (mm_interconnect_0_pwmonitor_i2c_avalon_slave_0_chipselect),       //                                           .chipselect
		.sysid_qsys_control_slave_address                 (mm_interconnect_0_sysid_qsys_control_slave_address),              //                   sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                (mm_interconnect_0_sysid_qsys_control_slave_readdata),             //                                           .readdata
		.timer_0_s1_address                               (mm_interconnect_0_timer_0_s1_address),                            //                                 timer_0_s1.address
		.timer_0_s1_write                                 (mm_interconnect_0_timer_0_s1_write),                              //                                           .write
		.timer_0_s1_readdata                              (mm_interconnect_0_timer_0_s1_readdata),                           //                                           .readdata
		.timer_0_s1_writedata                             (mm_interconnect_0_timer_0_s1_writedata),                          //                                           .writedata
		.timer_0_s1_chipselect                            (mm_interconnect_0_timer_0_s1_chipselect),                         //                                           .chipselect
		.uart_bt_avalon_rs232_slave_address               (mm_interconnect_0_uart_bt_avalon_rs232_slave_address),            //                 uart_bt_avalon_rs232_slave.address
		.uart_bt_avalon_rs232_slave_write                 (mm_interconnect_0_uart_bt_avalon_rs232_slave_write),              //                                           .write
		.uart_bt_avalon_rs232_slave_read                  (mm_interconnect_0_uart_bt_avalon_rs232_slave_read),               //                                           .read
		.uart_bt_avalon_rs232_slave_readdata              (mm_interconnect_0_uart_bt_avalon_rs232_slave_readdata),           //                                           .readdata
		.uart_bt_avalon_rs232_slave_writedata             (mm_interconnect_0_uart_bt_avalon_rs232_slave_writedata),          //                                           .writedata
		.uart_bt_avalon_rs232_slave_byteenable            (mm_interconnect_0_uart_bt_avalon_rs232_slave_byteenable),         //                                           .byteenable
		.uart_bt_avalon_rs232_slave_chipselect            (mm_interconnect_0_uart_bt_avalon_rs232_slave_chipselect)          //                                           .chipselect
	);

	Qsys_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                                   (clk_clk),                                                      //                                                 clk_0_clk.clk
		.mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_0_m0_address                           (mm_clock_crossing_bridge_0_m0_address),                        //                             mm_clock_crossing_bridge_0_m0.address
		.mm_clock_crossing_bridge_0_m0_waitrequest                       (mm_clock_crossing_bridge_0_m0_waitrequest),                    //                                                          .waitrequest
		.mm_clock_crossing_bridge_0_m0_burstcount                        (mm_clock_crossing_bridge_0_m0_burstcount),                     //                                                          .burstcount
		.mm_clock_crossing_bridge_0_m0_byteenable                        (mm_clock_crossing_bridge_0_m0_byteenable),                     //                                                          .byteenable
		.mm_clock_crossing_bridge_0_m0_read                              (mm_clock_crossing_bridge_0_m0_read),                           //                                                          .read
		.mm_clock_crossing_bridge_0_m0_readdata                          (mm_clock_crossing_bridge_0_m0_readdata),                       //                                                          .readdata
		.mm_clock_crossing_bridge_0_m0_readdatavalid                     (mm_clock_crossing_bridge_0_m0_readdatavalid),                  //                                                          .readdatavalid
		.mm_clock_crossing_bridge_0_m0_write                             (mm_clock_crossing_bridge_0_m0_write),                          //                                                          .write
		.mm_clock_crossing_bridge_0_m0_writedata                         (mm_clock_crossing_bridge_0_m0_writedata),                      //                                                          .writedata
		.mm_clock_crossing_bridge_0_m0_debugaccess                       (mm_clock_crossing_bridge_0_m0_debugaccess),                    //                                                          .debugaccess
		.LED_s1_address                                                  (mm_interconnect_1_led_s1_address),                             //                                                    LED_s1.address
		.LED_s1_write                                                    (mm_interconnect_1_led_s1_write),                               //                                                          .write
		.LED_s1_readdata                                                 (mm_interconnect_1_led_s1_readdata),                            //                                                          .readdata
		.LED_s1_writedata                                                (mm_interconnect_1_led_s1_writedata),                           //                                                          .writedata
		.LED_s1_chipselect                                               (mm_interconnect_1_led_s1_chipselect),                          //                                                          .chipselect
		.sonic_distance_0_avalon_slave_0_address                         (mm_interconnect_1_sonic_distance_0_avalon_slave_0_address),    //                           sonic_distance_0_avalon_slave_0.address
		.sonic_distance_0_avalon_slave_0_read                            (mm_interconnect_1_sonic_distance_0_avalon_slave_0_read),       //                                                          .read
		.sonic_distance_0_avalon_slave_0_readdata                        (mm_interconnect_1_sonic_distance_0_avalon_slave_0_readdata),   //                                                          .readdata
		.sonic_distance_0_avalon_slave_0_chipselect                      (mm_interconnect_1_sonic_distance_0_avalon_slave_0_chipselect)  //                                                          .chipselect
	);

	Qsys_irq_mapper irq_mapper (
		.clk           (pll_0_outclk0_clk),                  //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_0_outclk0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_0_outclk0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_0_outclk0_clk),                      //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk1_clk),                  //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
