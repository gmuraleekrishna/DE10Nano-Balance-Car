// Qsys_tb.v

// Generated using ACDS version 16.0 222

`timescale 1 ps / 1 ps
module Qsys_tb (
	);

	wire         qsys_inst_clk_bfm_clk_clk;                                              // Qsys_inst_clk_bfm:clk -> [Qsys_inst:clk_clk, Qsys_inst_reset_bfm:clk]
	wire   [0:0] qsys_inst_bts_tmd_connect_state_external_connection_bfm_conduit_export; // Qsys_inst_bts_tmd_connect_state_external_connection_bfm:sig_export -> Qsys_inst:bts_tmd_connect_state_external_connection_export
	wire         qsys_inst_buzzer_out_external_connection_export;                        // Qsys_inst:buzzer_out_external_connection_export -> Qsys_inst_buzzer_out_external_connection_bfm:sig_export
	wire   [1:0] qsys_inst_car_led_external_connection_export;                           // Qsys_inst:car_led_external_connection_export -> Qsys_inst_car_led_external_connection_bfm:sig_export
	wire  [11:0] qsys_inst_car_voltage_data_external_connection_bfm_conduit_export;      // Qsys_inst_car_voltage_data_external_connection_bfm:sig_export -> Qsys_inst:car_voltage_data_external_connection_export
	wire         qsys_inst_dc_motor_left_conduit_end_motor_p;                            // Qsys_inst:dc_motor_left_conduit_end_motor_p -> Qsys_inst_dc_motor_left_conduit_end_bfm:sig_motor_p
	wire         qsys_inst_dc_motor_left_conduit_end_motor_n;                            // Qsys_inst:dc_motor_left_conduit_end_motor_n -> Qsys_inst_dc_motor_left_conduit_end_bfm:sig_motor_n
	wire         qsys_inst_dc_motor_right_conduit_end_motor_p;                           // Qsys_inst:dc_motor_right_conduit_end_motor_p -> Qsys_inst_dc_motor_right_conduit_end_bfm:sig_motor_p
	wire         qsys_inst_dc_motor_right_conduit_end_motor_n;                           // Qsys_inst:dc_motor_right_conduit_end_motor_n -> Qsys_inst_dc_motor_right_conduit_end_bfm:sig_motor_n
	wire   [7:0] qsys_inst_led_external_connection_export;                               // Qsys_inst:led_external_connection_export -> Qsys_inst_led_external_connection_bfm:sig_export
	wire   [1:0] qsys_inst_motor_measure_left_conduit_end_bfm_conduit_ab;                // Qsys_inst_motor_measure_left_conduit_end_bfm:sig_ab -> Qsys_inst:motor_measure_left_conduit_end_ab
	wire   [1:0] qsys_inst_motor_measure_right_conduit_end_bfm_conduit_ab;               // Qsys_inst_motor_measure_right_conduit_end_bfm:sig_ab -> Qsys_inst:motor_measure_right_conduit_end_ab
	wire         qsys_inst_mpu_i2c_export_scl_pad_io;                                    // [] -> [Qsys_inst:mpu_i2c_export_scl_pad_io, Qsys_inst_mpu_i2c_export_bfm:sig_scl_pad_io]
	wire         qsys_inst_mpu_i2c_export_sda_pad_io;                                    // [] -> [Qsys_inst:mpu_i2c_export_sda_pad_io, Qsys_inst_mpu_i2c_export_bfm:sig_sda_pad_io]
	wire   [0:0] qsys_inst_mpu_int_external_connection_bfm_conduit_export;               // Qsys_inst_mpu_int_external_connection_bfm:sig_export -> Qsys_inst:mpu_int_external_connection_export
	wire   [0:0] qsys_inst_pmonitor_alert_external_connection_bfm_conduit_export;        // Qsys_inst_pmonitor_alert_external_connection_bfm:sig_export -> Qsys_inst:pmonitor_alert_external_connection_export
	wire         qsys_inst_pwmonitor_i2c_export_scl_pad_io;                              // [] -> [Qsys_inst:pwmonitor_i2c_export_scl_pad_io, Qsys_inst_pwmonitor_i2c_export_bfm:sig_scl_pad_io]
	wire         qsys_inst_pwmonitor_i2c_export_sda_pad_io;                              // [] -> [Qsys_inst:pwmonitor_i2c_export_sda_pad_io, Qsys_inst_pwmonitor_i2c_export_bfm:sig_sda_pad_io]
	wire   [0:0] qsys_inst_sonic_distance_0_conduit_end_bfm_conduit_echo;                // Qsys_inst_sonic_distance_0_conduit_end_bfm:sig_echo -> Qsys_inst:sonic_distance_0_conduit_end_echo
	wire         qsys_inst_sonic_distance_0_conduit_end_trigger;                         // Qsys_inst:sonic_distance_0_conduit_end_trigger -> Qsys_inst_sonic_distance_0_conduit_end_bfm:sig_trigger
	wire         qsys_inst_uart_bt_external_interface_txd;                               // Qsys_inst:uart_bt_external_interface_TXD -> Qsys_inst_uart_bt_external_interface_bfm:sig_TXD
	wire   [0:0] qsys_inst_uart_bt_external_interface_bfm_conduit_rxd;                   // Qsys_inst_uart_bt_external_interface_bfm:sig_RXD -> Qsys_inst:uart_bt_external_interface_RXD
	wire         qsys_inst_reset_bfm_reset_reset;                                        // Qsys_inst_reset_bfm:reset -> Qsys_inst:reset_reset_n

	Qsys qsys_inst (
		.bts_tmd_connect_state_external_connection_export (qsys_inst_bts_tmd_connect_state_external_connection_bfm_conduit_export), // bts_tmd_connect_state_external_connection.export
		.buzzer_out_external_connection_export            (qsys_inst_buzzer_out_external_connection_export),                        //            buzzer_out_external_connection.export
		.car_led_external_connection_export               (qsys_inst_car_led_external_connection_export),                           //               car_led_external_connection.export
		.car_voltage_data_external_connection_export      (qsys_inst_car_voltage_data_external_connection_bfm_conduit_export),      //      car_voltage_data_external_connection.export
		.clk_clk                                          (qsys_inst_clk_bfm_clk_clk),                                              //                                       clk.clk
		.dc_motor_left_conduit_end_motor_p                (qsys_inst_dc_motor_left_conduit_end_motor_p),                            //                 dc_motor_left_conduit_end.motor_p
		.dc_motor_left_conduit_end_motor_n                (qsys_inst_dc_motor_left_conduit_end_motor_n),                            //                                          .motor_n
		.dc_motor_right_conduit_end_motor_p               (qsys_inst_dc_motor_right_conduit_end_motor_p),                           //                dc_motor_right_conduit_end.motor_p
		.dc_motor_right_conduit_end_motor_n               (qsys_inst_dc_motor_right_conduit_end_motor_n),                           //                                          .motor_n
		.led_external_connection_export                   (qsys_inst_led_external_connection_export),                               //                   led_external_connection.export
		.motor_measure_left_conduit_end_ab                (qsys_inst_motor_measure_left_conduit_end_bfm_conduit_ab),                //            motor_measure_left_conduit_end.ab
		.motor_measure_right_conduit_end_ab               (qsys_inst_motor_measure_right_conduit_end_bfm_conduit_ab),               //           motor_measure_right_conduit_end.ab
		.mpu_i2c_export_scl_pad_io                        (qsys_inst_mpu_i2c_export_scl_pad_io),                                    //                            mpu_i2c_export.scl_pad_io
		.mpu_i2c_export_sda_pad_io                        (qsys_inst_mpu_i2c_export_sda_pad_io),                                    //                                          .sda_pad_io
		.mpu_int_external_connection_export               (qsys_inst_mpu_int_external_connection_bfm_conduit_export),               //               mpu_int_external_connection.export
		.pmonitor_alert_external_connection_export        (qsys_inst_pmonitor_alert_external_connection_bfm_conduit_export),        //        pmonitor_alert_external_connection.export
		.pwmonitor_i2c_export_scl_pad_io                  (qsys_inst_pwmonitor_i2c_export_scl_pad_io),                              //                      pwmonitor_i2c_export.scl_pad_io
		.pwmonitor_i2c_export_sda_pad_io                  (qsys_inst_pwmonitor_i2c_export_sda_pad_io),                              //                                          .sda_pad_io
		.reset_reset_n                                    (qsys_inst_reset_bfm_reset_reset),                                        //                                     reset.reset_n
		.sonic_distance_0_conduit_end_echo                (qsys_inst_sonic_distance_0_conduit_end_bfm_conduit_echo),                //              sonic_distance_0_conduit_end.echo
		.sonic_distance_0_conduit_end_trigger             (qsys_inst_sonic_distance_0_conduit_end_trigger),                         //                                          .trigger
		.uart_bt_external_interface_RXD                   (qsys_inst_uart_bt_external_interface_bfm_conduit_rxd),                   //                uart_bt_external_interface.RXD
		.uart_bt_external_interface_TXD                   (qsys_inst_uart_bt_external_interface_txd)                                //                                          .TXD
	);

	altera_conduit_bfm qsys_inst_bts_tmd_connect_state_external_connection_bfm (
		.sig_export (qsys_inst_bts_tmd_connect_state_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 qsys_inst_buzzer_out_external_connection_bfm (
		.sig_export (qsys_inst_buzzer_out_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm_0003 qsys_inst_car_led_external_connection_bfm (
		.sig_export (qsys_inst_car_led_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm_0004 qsys_inst_car_voltage_data_external_connection_bfm (
		.sig_export (qsys_inst_car_voltage_data_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) qsys_inst_clk_bfm (
		.clk (qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0005 qsys_inst_dc_motor_left_conduit_end_bfm (
		.sig_motor_p (qsys_inst_dc_motor_left_conduit_end_motor_p), // conduit.motor_p
		.sig_motor_n (qsys_inst_dc_motor_left_conduit_end_motor_n)  //        .motor_n
	);

	altera_conduit_bfm_0005 qsys_inst_dc_motor_right_conduit_end_bfm (
		.sig_motor_p (qsys_inst_dc_motor_right_conduit_end_motor_p), // conduit.motor_p
		.sig_motor_n (qsys_inst_dc_motor_right_conduit_end_motor_n)  //        .motor_n
	);

	altera_conduit_bfm_0006 qsys_inst_led_external_connection_bfm (
		.sig_export (qsys_inst_led_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm_0007 qsys_inst_motor_measure_left_conduit_end_bfm (
		.sig_ab (qsys_inst_motor_measure_left_conduit_end_bfm_conduit_ab)  // conduit.ab
	);

	altera_conduit_bfm_0007 qsys_inst_motor_measure_right_conduit_end_bfm (
		.sig_ab (qsys_inst_motor_measure_right_conduit_end_bfm_conduit_ab)  // conduit.ab
	);

	altera_conduit_bfm_0008 qsys_inst_mpu_i2c_export_bfm (
		.sig_scl_pad_io (qsys_inst_mpu_i2c_export_scl_pad_io), // conduit.scl_pad_io
		.sig_sda_pad_io (qsys_inst_mpu_i2c_export_sda_pad_io)  //        .sda_pad_io
	);

	altera_conduit_bfm qsys_inst_mpu_int_external_connection_bfm (
		.sig_export (qsys_inst_mpu_int_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm qsys_inst_pmonitor_alert_external_connection_bfm (
		.sig_export (qsys_inst_pmonitor_alert_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0008 qsys_inst_pwmonitor_i2c_export_bfm (
		.sig_scl_pad_io (qsys_inst_pwmonitor_i2c_export_scl_pad_io), // conduit.scl_pad_io
		.sig_sda_pad_io (qsys_inst_pwmonitor_i2c_export_sda_pad_io)  //        .sda_pad_io
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) qsys_inst_reset_bfm (
		.reset (qsys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (qsys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0009 qsys_inst_sonic_distance_0_conduit_end_bfm (
		.sig_echo    (qsys_inst_sonic_distance_0_conduit_end_bfm_conduit_echo), // conduit.echo
		.sig_trigger (qsys_inst_sonic_distance_0_conduit_end_trigger)           //        .trigger
	);

	altera_conduit_bfm_0010 qsys_inst_uart_bt_external_interface_bfm (
		.sig_RXD (qsys_inst_uart_bt_external_interface_bfm_conduit_rxd), // conduit.RXD
		.sig_TXD (qsys_inst_uart_bt_external_interface_txd)              //        .TXD
	);

endmodule
