// (C) 2001-2016 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// $Id: //acds/main/ip/sopc/components/verification/altera_tristate_conduit_bfm/altera_tristate_conduit_bfm.sv.terp#7 $
// $Revision: #7 $
// $Date: 2010/08/05 $
// $Author: klong $
//-----------------------------------------------------------------------------
// =head1 NAME
// altera_conduit_bfm
// =head1 SYNOPSIS
// Bus Functional Model (BFM) for a Standard Conduit BFM
//-----------------------------------------------------------------------------
// =head1 DESCRIPTION
// This is a Bus Functional Model (BFM) for a Standard Conduit Master.
// This BFM sampled the input/bidirection port value or driving user's value to 
// output ports when user call the API.  
// This BFM's HDL is been generated through terp file in Qsys/SOPC Builder.
// Generation parameters:
// output_name:                                       altera_conduit_bfm_0009
// role:width:direction:                              echo:1:output,trigger:1:input
// 0
//-----------------------------------------------------------------------------
`timescale 1 ps / 1 ps

module altera_conduit_bfm_0009
(
   sig_echo,
   sig_trigger
);

   //--------------------------------------------------------------------------
   // =head1 PINS 
   // =head2 User defined interface
   //--------------------------------------------------------------------------
   output sig_echo;
   input sig_trigger;

   // synthesis translate_off
   import verbosity_pkg::*;
   
   typedef logic ROLE_echo_t;
   typedef logic ROLE_trigger_t;

   reg sig_echo_temp;
   reg sig_echo_out;
   logic [0 : 0] sig_trigger_in;
   logic [0 : 0] sig_trigger_local;

   //--------------------------------------------------------------------------
   // =head1 Public Methods API
   // =pod
   // This section describes the public methods in the application programming
   // interface (API). The application program interface provides methods for 
   // a testbench which instantiates, controls and queries state in this BFM 
   // component. Test programs must only use these public access methods and 
   // events to communicate with this BFM component. The API and module pins
   // are the only interfaces of this component that are guaranteed to be
   // stable. The API will be maintained for the life of the product. 
   // While we cannot prevent a test program from directly accessing internal
   // tasks, functions, or data private to the BFM, there is no guarantee that
   // these will be present in the future. In fact, it is best for the user
   // to assume that the underlying implementation of this component can 
   // and will change.
   // =cut
   //--------------------------------------------------------------------------
   
   event signal_input_trigger_change;
   
   function automatic string get_version();  // public
      // Return BFM version string. For example, version 9.1 sp1 is "9.1sp1" 
      string ret_version = "16.0";
      return ret_version;
   endfunction

   // -------------------------------------------------------
   // echo
   // -------------------------------------------------------

   function automatic void set_echo (
      ROLE_echo_t new_value
   );
      // Drive the new value to echo.
      
      $sformat(message, "%m: method called arg0 %0d", new_value); 
      print(VERBOSITY_DEBUG, message);
      
      sig_echo_temp = new_value;
   endfunction

   // -------------------------------------------------------
   // trigger
   // -------------------------------------------------------
   function automatic ROLE_trigger_t get_trigger();
   
      // Gets the trigger input value.
      $sformat(message, "%m: called get_trigger");
      print(VERBOSITY_DEBUG, message);
      return sig_trigger_in;
      
   endfunction

   assign sig_echo = sig_echo_temp;
   assign sig_trigger_in = sig_trigger;


   always @(sig_trigger_in) begin
      if (sig_trigger_local != sig_trigger_in)
         -> signal_input_trigger_change;
      sig_trigger_local = sig_trigger_in;
   end
   


// synthesis translate_on

endmodule

